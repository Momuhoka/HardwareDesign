//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Thu Jun 13 09:45:30 2024

module music_SP (dout, clk, oce, ce, reset, wre, ad, din);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [11:0] ad;
input [15:0] din;

wire [27:0] sp_inst_0_dout_w;
wire [27:0] sp_inst_1_dout_w;
wire [27:0] sp_inst_2_dout_w;
wire [27:0] sp_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 4;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hB082780488270F41F088A8F08717A4AA0FA8AB8F188A8F488FF47B100FBFAFAF;
defparam sp_inst_0.INIT_RAM_01 = 256'hA178B4F18B178F0FB8780B24F2FF0F207288F8F208F08B87017F82112F84171F;
defparam sp_inst_0.INIT_RAM_02 = 256'hF87AAA88F14F77874448B41FF088ABF80F2808F42A7F04AFF78F7BFF0011182F;
defparam sp_inst_0.INIT_RAM_03 = 256'h1784FFB8181882F7A4F8A77848AB44B844F242A8428BA782AFB0B27A8BF8027A;
defparam sp_inst_0.INIT_RAM_04 = 256'h7071AF88B778228F77488FF2718A144F7272F2410BFA7F12F728AF8B24F440FF;
defparam sp_inst_0.INIT_RAM_05 = 256'h41B4A17B42FA21224882FF7A2F1B1AFA880FA210220A4F4F822178F78A77F17B;
defparam sp_inst_0.INIT_RAM_06 = 256'h04B242A08072AFF8B8F0A7FF41B8781AF4014A8A7878BAAFA27F08FF4AFF2AF0;
defparam sp_inst_0.INIT_RAM_07 = 256'hF88A07820810B81FA24B0014F878412A2A88A8F1288F7880BFBBF08A8FAF82A7;
defparam sp_inst_0.INIT_RAM_08 = 256'h081744217F2F1AF7148BA08AB0AF7BFAF10FB020FBBF7FF1FA7487800B040AF0;
defparam sp_inst_0.INIT_RAM_09 = 256'hB7F87201F48ABBA801880112AFFF14F71274882B218AF728FFA4F2A727F278BF;
defparam sp_inst_0.INIT_RAM_0A = 256'h87F14F1B8888A7FA40FBB10B08BF8B407788280A2478F17BFF8080F8FF77AF8F;
defparam sp_inst_0.INIT_RAM_0B = 256'h8887FFB24022A0B81F21B22A847A778AFB88AB08F7FBFAF788B4F741480FFAF4;
defparam sp_inst_0.INIT_RAM_0C = 256'h7187888828274AA87BFA00A148F178F81AB021F4B87FFBF4A1FA74078B488118;
defparam sp_inst_0.INIT_RAM_0D = 256'h401AF7A88248AB70AB81780F80FA787F7B2482F08F1B840B28F2748B7AF0F877;
defparam sp_inst_0.INIT_RAM_0E = 256'hB7A0F1A2A1887247140A8181AB87871B211A4FF2124874B20A2FBF848F721728;
defparam sp_inst_0.INIT_RAM_0F = 256'h804481FAF42A7204A010FFA04F7BBFF281148B8BBAB77A21287A47A8B71F8A2F;
defparam sp_inst_0.INIT_RAM_10 = 256'h7F0BF2288A2871027A887A1088F0A0B424BBFF441F888818784BABFF8BF71807;
defparam sp_inst_0.INIT_RAM_11 = 256'h24A10417BB80F127ABA072878278B17F74172878A011F78FB2F8AFAF471AFF28;
defparam sp_inst_0.INIT_RAM_12 = 256'hFF77F70BFFBA7F8FAF0B07F7488F2F8724200821FFAF888BF280A8AF02AB78B4;
defparam sp_inst_0.INIT_RAM_13 = 256'h427BA2B48FB7784BAF0FF0F48B04880488A88011210F2142182F01F1B881F71F;
defparam sp_inst_0.INIT_RAM_14 = 256'h144FAB41B24F1B2712218041F8708800FA844BF8F08244F8F1122FF1288784A8;
defparam sp_inst_0.INIT_RAM_15 = 256'h1428FA0BFB4FFF8287B207B8BF777810F20AF000144BA101B1FA400B8BFAFF27;
defparam sp_inst_0.INIT_RAM_16 = 256'h87817270B708F08F0712F84F77070B128BFF820FA007FA2FF4A08010047FF447;
defparam sp_inst_0.INIT_RAM_17 = 256'hFA8A1444F4F80F412AB24A244272B2A0B8F2828A2BFFA4442BF7401B7A248AB7;
defparam sp_inst_0.INIT_RAM_18 = 256'h8888B7222488B148444AA028F8F024FBA241F44BF2111AAF2BFAA081F7411178;
defparam sp_inst_0.INIT_RAM_19 = 256'h10444BBFF882FAFAFAF77144BF1F0F171FAA274AAA1B0A817AA7F28FFFA47BB4;
defparam sp_inst_0.INIT_RAM_1A = 256'h0B2F4B47F8A8FF88AA8FA0B8FA42177F8BA0F48F2A24AA1781870FABFA218F4A;
defparam sp_inst_0.INIT_RAM_1B = 256'h844B188F8A84A28F4F4777FF48882012A0B0FAB10BFA1A841721A082B4F80F7B;
defparam sp_inst_0.INIT_RAM_1C = 256'h7A878101A7FA11880B2F8B77FAA7FAFAF08784B888811FBF88BFF7A2F7808227;
defparam sp_inst_0.INIT_RAM_1D = 256'h887A88FFF0A8F247278FF808B8FB01748804FA08F8A7FFF4F8B184F2F401F784;
defparam sp_inst_0.INIT_RAM_1E = 256'hFF172F884AF8871828A84821870842424801812F4FA8FFFA880F0087042FF8AA;
defparam sp_inst_0.INIT_RAM_1F = 256'h82B24F842BA2B84A8FFAB871884248220A7F082F8A1AB7728F082110818F4888;
defparam sp_inst_0.INIT_RAM_20 = 256'h2F221F0BA04F0B2AA8724F2008248B1104288A7FF171202F708A8F80AFFF821A;
defparam sp_inst_0.INIT_RAM_21 = 256'h0782F111A8747882B011BBA8082181828AB880448AF8A28B8F82BF47AFFF8108;
defparam sp_inst_0.INIT_RAM_22 = 256'hF2A74A8704BF7F4A2FF4FB427FFFF478F0AFBF7B0F8F218B27B0AA4BBA18F4F1;
defparam sp_inst_0.INIT_RAM_23 = 256'h028BFF82024022A74B1278121FAF128FF728F8A1412F1F8170FAFF7244FFB2A4;
defparam sp_inst_0.INIT_RAM_24 = 256'h0A2018A180700880F187AFFFF10B0808BFF2F14A708F4B84AA4AB18A4F8FF817;
defparam sp_inst_0.INIT_RAM_25 = 256'h8B188A4288288F4F8FA80F4228F0F848B01BBF8F8F2088FA10418F8A77447117;
defparam sp_inst_0.INIT_RAM_26 = 256'hF0872488048F8BFF0871278A1A488201A84282B2FF2A40BAB8F1F81A81278FA0;
defparam sp_inst_0.INIT_RAM_27 = 256'hFFF88A04B02B800B17142F28F28810A808710F80A1F2BA2441AFB8A7AAB02811;
defparam sp_inst_0.INIT_RAM_28 = 256'h742A88FF0A20FF7FB20720FF4401B1F4FB22B08BB08A0F7FF78F84F72A7B1B00;
defparam sp_inst_0.INIT_RAM_29 = 256'h01BA82AFF2FFB08F1F72A4AB8A87AF80F87F84AF48B18BBF1202B0F102887AB4;
defparam sp_inst_0.INIT_RAM_2A = 256'h84BB047208B8B1F0A01021FB14A8BFABF7BA12F72FF4A8128F80FA11FFB717BB;
defparam sp_inst_0.INIT_RAM_2B = 256'h7217740F887884AFF410F874A087782FBBF4FFF81B72B1701AF8F8B0884FF14A;
defparam sp_inst_0.INIT_RAM_2C = 256'h4401AA2147AF282A877F4A7F81F1F2A11FF7408780B820A8F044B4AAFF7FA81A;
defparam sp_inst_0.INIT_RAM_2D = 256'h07F8F0B4B21A18F4174A87B84FA8F8028847A040B1F410B7F87480AF82AF7228;
defparam sp_inst_0.INIT_RAM_2E = 256'h8FF0BB820BB188FF8781228FABAB78740B8FFF0A14108017028B1002471F80FF;
defparam sp_inst_0.INIT_RAM_2F = 256'hBA4028708A04841808A4FFA7FB478FBFFA712FF2F78AF48F8F8B8F84F8102A27;
defparam sp_inst_0.INIT_RAM_30 = 256'h4A48AFF8178FA7F7B2F08888F8ABF888A1824F47717B4FBB42F7FAF887F2B727;
defparam sp_inst_0.INIT_RAM_31 = 256'h0084B847F27001F12F8B24AA028F784FB18F1818AFF102F8884A80A7B0F8F2B8;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 4;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h6877898B997888BAB899A78898A8ABAA88A7A69BA97A9BB97B8B86A88868ABAB;
defparam sp_inst_1.INIT_RAM_01 = 256'hAA876BBA76A878886787867B87BB8B788779B98787B896988A8B77AA787BA8AB;
defparam sp_inst_1.INIT_RAM_02 = 256'h898AAA77BABB8898BBB76BAB8899A6B7887987BB7A8B8BAB8878868888AAA97B;
defparam sp_inst_1.INIT_RAM_03 = 256'hA87BBB69A9A77788AB87A887B7A6BB67BBB7B7A7B796A897AB68678A96B9878A;
defparam sp_inst_1.INIT_RAM_04 = 256'h888AA8796887777888B77BB78A7AABB8878787BA86BA88A78879AB967BBBB888;
defparam sp_inst_1.INIT_RAM_05 = 256'hBA6BAA86B7BA7A77B977B88A78A6AABA778BA7A8778ABBBB777A89B87A888A86;
defparam sp_inst_1.INIT_RAM_06 = 256'h8B67B7A87887A88767B8A8B8BA6789AA8B8ABA7A87896AABA78B87B8BA8B7AB8;
defparam sp_inst_1.INIT_RAM_07 = 256'h879A889789A869ABA7B688AB8789BA7A7A77A7BA799B89786866889A9BAB77A8;
defparam sp_inst_1.INIT_RAM_08 = 256'h89A8BB7A887BAAB8AB96A87A68AB868ABA886878B66B8B8ABA8B9878868B8AB8;
defparam sp_inst_1.INIT_RAM_09 = 256'h6887878A8B9A66A98A778AA7AB88ABB8A78B99767A7A8877BBAB87A878B78968;
defparam sp_inst_1.INIT_RAM_0A = 256'h988ABBA69979A88AB8866A86876B96B88899778A7B87BA868B7878898888AB98;
defparam sp_inst_1.INIT_RAM_0B = 256'h9798B867B877A869AB7A677A7B8A887AB679A687B8868AB8796BB8BAB98B8A8B;
defparam sp_inst_1.INIT_RAM_0C = 256'h8A7877997778BAA786BA88AAB98A87B7AA687ABB698B86BBAA8A8B8876B99AA9;
defparam sp_inst_1.INIT_RAM_0D = 256'hB8AA88A977B7A688A67A878B988A8988867B77B89BA67B8677B78B968A888788;
defparam sp_inst_1.INIT_RAM_0E = 256'h68A8BAA7AA7787B8AB8A7A9AA69878A67AAAB8B7A7B98B678A7B6B9B9887A879;
defparam sp_inst_1.INIT_RAM_0F = 256'h98BB9ABA8B7A878BA8A8BBA8B88668877AAB96966A688A7A798AB8A768AB7A78;
defparam sp_inst_1.INIT_RAM_10 = 256'h8B86B7799A798A878A798AA899B8A86B7B6688BBA87777A787B6A68B76B8A988;
defparam sp_inst_1.INIT_RAM_11 = 256'h7BAA8BA86678BA78A6A8877877896A888BA87987A8AAB87867B7ABA8B8AABB77;
defparam sp_inst_1.INIT_RAM_12 = 256'hBB88B8868B6A8B9BAB8688B8B79B78987B78877ABBA899768778A9AB87A6896B;
defparam sp_inst_1.INIT_RAM_13 = 256'hB786A76B7B6889B6AB8888BB968B978B97A778AA7A8B7AB7A7788ABA679AB8A8;
defparam sp_inst_1.INIT_RAM_14 = 256'hABB8A6BA67B8A678A77A98BA89889988BA9BB6B98877BBB78AA7788A77987BA7;
defparam sp_inst_1.INIT_RAM_15 = 256'hAB798A86B6B88B9798678867688887A8B78A8888ABB6AA8A6ABAB88696BAB878;
defparam sp_inst_1.INIT_RAM_16 = 256'h789A87886887887888A7B7B8888886A79688978BA8888A7BBBA878A88B8BBBB8;
defparam sp_inst_1.INIT_RAM_17 = 256'hBA9AABBBBBB788BA7A67BA7BB78767A867B7779A76BBABBB7688B8A68A7B9A68;
defparam sp_inst_1.INIT_RAM_18 = 256'h777968777B976AB7BBBAA87789B87BB6A7BABBB6B7AAAAAB768AA87AB8BAAA89;
defparam sp_inst_1.INIT_RAM_19 = 256'hA8BBB66B89978A8A8A888ABB68A88BA8A8AA78BAAAA68A7A8AA88778B8AB866B;
defparam sp_inst_1.INIT_RAM_1A = 256'h8678B6B889A9B877AA9BA869BAB7A88B76A88B787A7BAAA87A988BA68A7A98BA;
defparam sp_inst_1.INIT_RAM_1B = 256'h7BB6A99B7A7BA798BBB88888B79778A7A868BA6A86BAAA9BA87AA8976BB98886;
defparam sp_inst_1.INIT_RAM_1C = 256'h8A789A8AA88AAA97867B9688BAA88A8A88987B67779AAB68796888A788787778;
defparam sp_inst_1.INIT_RAM_1D = 256'h998A99B888A9B7B87898B78767868A8B798BBA8989A888BB876A9BB7BB8AB87B;
defparam sp_inst_1.INIT_RAM_1E = 256'h88A87B99BA8778A977A9B97A7889B7B7B98A9A78BBA988BA978B88788B7BB7AA;
defparam sp_inst_1.INIT_RAM_1F = 256'h7767BB9B76A769BA98BA698A79B7B9778A8B89787AAA68879B897AA87A9BB777;
defparam sp_inst_1.INIT_RAM_20 = 256'h7877A886A8BB867AA787BB78877B96AA8B799A8BBA8A7878889A9B78ABB897AA;
defparam sp_inst_1.INIT_RAM_21 = 256'h88978AAAA78B879768AA66A7897A7A777A6778BB9A87A796787768B8AB889A89;
defparam sp_inst_1.INIT_RAM_22 = 256'hB7A8BA988B6B8BBA788B86B788BBBB87B8AB688688987A767868AAB66AA9BBBA;
defparam sp_inst_1.INIT_RAM_23 = 256'h8796B87787B877A8B6A787A7ABA8A79BB87787AABA78A89A888AB887BBB867AB;
defparam sp_inst_1.INIT_RAM_24 = 256'h8A78A9AA988889988A98AB8BBA8689896B878ABA8898B69BAABA6A9ABB7B87A8;
defparam sp_inst_1.INIT_RAM_25 = 256'h76A77AB779777BB89BA78BB777B887B968A66B789B78978AA8BA789A88BB8AA8;
defparam sp_inst_1.INIT_RAM_26 = 256'h88787B798B987688878A789AAAB9778AA7B77767887AB86A698A87AA9A789BA8;
defparam sp_inst_1.INIT_RAM_27 = 256'h8B899A8B68767886A8AB7B798797A8A9898A8898AAB76A7BBAA867A8AA6879AA;
defparam sp_inst_1.INIT_RAM_28 = 256'h8B7A97888A78888867887888BB8A6ABB86776896687A888BB8787B887A86A688;
defparam sp_inst_1.INIT_RAM_29 = 256'h8A6A97AB87B86878A887ABA67A98A878B98B7BA8B96A7668A78768BA87798A6B;
defparam sp_inst_1.INIT_RAM_2A = 256'h7B668B8787696AB8A8A87AB6ABA968A6886AA78878BBA9A77B78BAAAB868A866;
defparam sp_inst_1.INIT_RAM_2B = 256'h87A88B8879899BABBBA8878BA878877B668B8B87A6876A88AA89876897BBBABA;
defparam sp_inst_1.INIT_RAM_2C = 256'hBB8AAA7AB8AB777A988BBA8B9A8AB7AAA8B8B878786978A788BB6BAABB88A9AA;
defparam sp_inst_1.INIT_RAM_2D = 256'h88B9886B67AAA98BA8BA7869BBA9B98777B8A8B86A8BA868898B78A897A88779;
defparam sp_inst_1.INIT_RAM_2E = 256'h98B86677866A778B989A779BA6A6878B869BB88AABA898A88776A887B8A878BB;
defparam sp_inst_1.INIT_RAM_2F = 256'h6AB877889A8B7BA987AB88A8B6B89B68BA8A7BB7889A8B7B9876987BB7A87A78;
defparam sp_inst_1.INIT_RAM_30 = 256'hBAB9A889A878A88867B87999B7A68977AA97B8B88A86BB66B7B88AB798B76878;
defparam sp_inst_1.INIT_RAM_31 = 256'h009B67B887888A8A78967BAA879B89B86A78A7A9AB8A87B797BA98A868B98767;
defparam sp_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:8]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 4;
defparam sp_inst_2.BLK_SEL = 3'b000;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[27:0],dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:12]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 4;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //music_SP
