module gw_gao(
    \speaker_music/addr[6] ,
    \speaker_music/addr[5] ,
    \speaker_music/addr[4] ,
    \speaker_music/addr[3] ,
    \speaker_music/addr[2] ,
    \speaker_music/addr[1] ,
    \speaker_music/addr[0] ,
    \speaker_music/data[15] ,
    \speaker_music/data[14] ,
    \speaker_music/data[13] ,
    \speaker_music/data[12] ,
    \speaker_music/data[11] ,
    \speaker_music/data[10] ,
    \speaker_music/data[9] ,
    \speaker_music/data[8] ,
    \speaker_music/data[7] ,
    \speaker_music/data[6] ,
    \speaker_music/data[5] ,
    \speaker_music/data[4] ,
    \speaker_music/data[3] ,
    \speaker_music/data[2] ,
    \speaker_music/data[1] ,
    \speaker_music/data[0] ,
    sys_clk,
    sys_rst_n,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \speaker_music/addr[6] ;
input \speaker_music/addr[5] ;
input \speaker_music/addr[4] ;
input \speaker_music/addr[3] ;
input \speaker_music/addr[2] ;
input \speaker_music/addr[1] ;
input \speaker_music/addr[0] ;
input \speaker_music/data[15] ;
input \speaker_music/data[14] ;
input \speaker_music/data[13] ;
input \speaker_music/data[12] ;
input \speaker_music/data[11] ;
input \speaker_music/data[10] ;
input \speaker_music/data[9] ;
input \speaker_music/data[8] ;
input \speaker_music/data[7] ;
input \speaker_music/data[6] ;
input \speaker_music/data[5] ;
input \speaker_music/data[4] ;
input \speaker_music/data[3] ;
input \speaker_music/data[2] ;
input \speaker_music/data[1] ;
input \speaker_music/data[0] ;
input sys_clk;
input sys_rst_n;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \speaker_music/addr[6] ;
wire \speaker_music/addr[5] ;
wire \speaker_music/addr[4] ;
wire \speaker_music/addr[3] ;
wire \speaker_music/addr[2] ;
wire \speaker_music/addr[1] ;
wire \speaker_music/addr[0] ;
wire \speaker_music/data[15] ;
wire \speaker_music/data[14] ;
wire \speaker_music/data[13] ;
wire \speaker_music/data[12] ;
wire \speaker_music/data[11] ;
wire \speaker_music/data[10] ;
wire \speaker_music/data[9] ;
wire \speaker_music/data[8] ;
wire \speaker_music/data[7] ;
wire \speaker_music/data[6] ;
wire \speaker_music/data[5] ;
wire \speaker_music/data[4] ;
wire \speaker_music/data[3] ;
wire \speaker_music/data[2] ;
wire \speaker_music/data[1] ;
wire \speaker_music/data[0] ;
wire sys_clk;
wire sys_rst_n;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\speaker_music/addr[6] ,\speaker_music/addr[5] ,\speaker_music/addr[4] ,\speaker_music/addr[3] ,\speaker_music/addr[2] ,\speaker_music/addr[1] ,\speaker_music/addr[0] }),
    .data_i({\speaker_music/addr[6] ,\speaker_music/addr[5] ,\speaker_music/addr[4] ,\speaker_music/addr[3] ,\speaker_music/addr[2] ,\speaker_music/addr[1] ,\speaker_music/addr[0] ,\speaker_music/data[15] ,\speaker_music/data[14] ,\speaker_music/data[13] ,\speaker_music/data[12] ,\speaker_music/data[11] ,\speaker_music/data[10] ,\speaker_music/data[9] ,\speaker_music/data[8] ,\speaker_music/data[7] ,\speaker_music/data[6] ,\speaker_music/data[5] ,\speaker_music/data[4] ,\speaker_music/data[3] ,\speaker_music/data[2] ,\speaker_music/data[1] ,\speaker_music/data[0] ,sys_clk,sys_rst_n}),
    .clk_i(sys_clk)
);

endmodule
